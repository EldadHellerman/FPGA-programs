module main(input clk, [1:0] buttons, output reg [5:0] leds);

endmodule
